package dma_ral_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "intr.sv"
	`include "ctrl.sv"
	`include "io_addr.sv"
	`include "mem_addr.sv"
	
	`include "dma_reg_model.sv"
endpackage